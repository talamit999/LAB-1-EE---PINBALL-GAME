module BlockBitMap (

					input	logic	clk, 
					input	logic	resetN, 
					input logic	[10:0] pixelX,// offset from top left  position 
					input logic	[10:0] pixelY, 
					input logic [3:0] level, // current level 
 
					output	logic	[7:0] RGBout  //rgb value from the bitmap 
 ) ; 
 
 
// generating the bitmap 

 

localparam logic [7:0] TRANSPARENT_ENCODING = 8'h00 ;// RGB value in the bitmap representing a transparent pixel  
logic[0:31][0:31][7:0] object_colors = {
	{8'hc0,8'h40,8'h80,8'h40,8'h40,8'h80,8'h40,8'h40,8'hc0,8'h40,8'h80,8'hc0,8'h40,8'h80,8'h80,8'h40,8'hc0,8'h40,8'h40,8'hc0,8'h00,8'h80,8'hc0,8'h40,8'h80,8'h40,8'h40,8'hc0,8'h00,8'h80,8'hc0,8'h40},
	{8'h80,8'hc0,8'h40,8'h80,8'h40,8'h40,8'hc0,8'h40,8'h40,8'hc0,8'h40,8'h80,8'hc0,8'h40,8'h80,8'h80,8'h40,8'hc0,8'h00,8'h40,8'hc0,8'h00,8'h80,8'hc0,8'h40,8'hc0,8'h40,8'h40,8'hc0,8'h40,8'h80,8'h80},
	{8'h40,8'h80,8'hc0,8'h40,8'h80,8'h40,8'h40,8'hc0,8'h40,8'h40,8'hc0,8'h00,8'h80,8'hc0,8'h40,8'h80,8'h80,8'h40,8'hc0,8'h00,8'h40,8'hc0,8'h00,8'h80,8'h80,8'h40,8'hc0,8'h40,8'h40,8'hc0,8'h40,8'h80},
	{8'hc0,8'h40,8'h80,8'hc0,8'h40,8'h80,8'h40,8'h40,8'hc0,8'h40,8'h40,8'hc0,8'h40,8'h80,8'hc0,8'h40,8'h80,8'h40,8'h40,8'hc0,8'h00,8'h80,8'hc0,8'h40,8'h80,8'h80,8'h40,8'hc0,8'h40,8'h40,8'hc0,8'h40},
	{8'h80,8'hc0,8'h40,8'h80,8'hc0,8'h40,8'hc0,8'h40,8'h40,8'hc0,8'h00,8'h80,8'hc0,8'h40,8'h80,8'hc0,8'h40,8'h80,8'h40,8'h40,8'hc0,8'h00,8'h80,8'hc0,8'h40,8'h80,8'h80,8'h40,8'hc0,8'h00,8'h40,8'hc0},
	{8'h40,8'h80,8'hc0,8'h40,8'h80,8'hc0,8'h40,8'hc0,8'h00,8'h40,8'hc0,8'h00,8'h80,8'hc0,8'h40,8'h80,8'hc0,8'h40,8'hc0,8'h40,8'h40,8'hc0,8'h00,8'h80,8'hc0,8'h40,8'h80,8'h40,8'h40,8'hc0,8'h40,8'h40},
	{8'hc0,8'h40,8'h80,8'hc0,8'h40,8'h80,8'hc0,8'h40,8'hc0,8'h40,8'h80,8'hc0,8'h40,8'h80,8'hc0,8'h40,8'h80,8'hc0,8'h40,8'h80,8'h40,8'h40,8'hc0,8'h00,8'h80,8'hc0,8'h40,8'hc0,8'h40,8'h40,8'hc0,8'h00},
	{8'h80,8'hc0,8'h40,8'h80,8'hc0,8'h40,8'h80,8'hc0,8'h40,8'hc0,8'h40,8'h80,8'hc0,8'h00,8'h80,8'hc0,8'h40,8'h80,8'hc0,8'h40,8'hc0,8'h40,8'h40,8'hc0,8'h40,8'h80,8'hc0,8'h40,8'hc0,8'h40,8'h80,8'hc0},
	{8'h00,8'h80,8'hc0,8'h40,8'h80,8'hc0,8'h40,8'h80,8'hc0,8'h40,8'hc0,8'h40,8'h80,8'hc0,8'h40,8'h80,8'hc0,8'h40,8'h80,8'hc0,8'h40,8'hc0,8'h40,8'h40,8'hc0,8'h40,8'h80,8'hc0,8'h40,8'hc0,8'h00,8'h80},
	{8'hc0,8'h40,8'h80,8'hc0,8'h00,8'h80,8'hc0,8'h40,8'h80,8'hc0,8'h40,8'hc0,8'h00,8'h80,8'hc0,8'h40,8'h80,8'hc0,8'h40,8'h80,8'hc0,8'h40,8'hc0,8'h00,8'h80,8'hc0,8'h40,8'h80,8'h80,8'h40,8'hc0,8'h00},
	{8'h80,8'hc0,8'h00,8'h80,8'hc0,8'h00,8'h80,8'hc0,8'h40,8'h80,8'hc0,8'h40,8'hc0,8'h00,8'h80,8'hc0,8'h40,8'h80,8'hc0,8'h40,8'h80,8'hc0,8'h40,8'hc0,8'h40,8'h80,8'hc0,8'h40,8'h80,8'hc0,8'h40,8'hc0},
	{8'h40,8'h80,8'hc0,8'h40,8'h80,8'hc0,8'h40,8'h80,8'hc0,8'h40,8'h80,8'h80,8'h40,8'hc0,8'h40,8'h80,8'hc0,8'h40,8'h80,8'hc0,8'h40,8'h80,8'hc0,8'h40,8'hc0,8'h00,8'h80,8'hc0,8'h40,8'h80,8'h80,8'h40},
	{8'hc0,8'h40,8'h80,8'hc0,8'h40,8'h80,8'hc0,8'h40,8'h80,8'hc0,8'h40,8'h80,8'h80,8'h40,8'hc0,8'h40,8'h80,8'hc0,8'h40,8'h80,8'hc0,8'h40,8'hc0,8'hc0,8'h40,8'hc0,8'h00,8'h80,8'hc0,8'h40,8'hc0,8'h80},
	{8'h40,8'hc0,8'h00,8'h80,8'hc0,8'h00,8'h80,8'hc0,8'h40,8'h80,8'hc0,8'h40,8'hc0,8'h80,8'h40,8'hc0,8'h00,8'h80,8'hc0,8'h40,8'h80,8'h80,8'h40,8'hc0,8'h80,8'h40,8'hc0,8'h00,8'h80,8'hc0,8'h40,8'hc0},
	{8'h80,8'h40,8'hc0,8'h00,8'h80,8'hc0,8'h40,8'h80,8'hc0,8'h40,8'h80,8'hc0,8'h40,8'h80,8'h80,8'h40,8'hc0,8'h00,8'h80,8'hc0,8'h40,8'h80,8'h80,8'h40,8'hc0,8'h80,8'h40,8'hc0,8'h40,8'h80,8'hc0,8'h40},
	{8'hc0,8'h80,8'h40,8'hc0,8'h00,8'h80,8'hc0,8'h40,8'h80,8'hc0,8'h40,8'h80,8'h80,8'h40,8'hc0,8'h80,8'h40,8'hc0,8'h40,8'h80,8'hc0,8'h40,8'h80,8'h80,8'h40,8'hc0,8'h40,8'h40,8'hc0,8'h40,8'h80,8'hc0},
	{8'h40,8'hc0,8'h80,8'h40,8'hc0,8'h40,8'h80,8'hc0,8'h40,8'h80,8'hc0,8'h40,8'h80,8'hc0,8'h40,8'h80,8'h80,8'h40,8'hc0,8'h40,8'h80,8'hc0,8'h40,8'h80,8'h80,8'h40,8'hc0,8'h80,8'h40,8'hc0,8'h40,8'h80},
	{8'hc0,8'h40,8'hc0,8'h80,8'h40,8'hc0,8'h40,8'h80,8'hc0,8'h40,8'h80,8'hc0,8'h40,8'h80,8'hc0,8'h40,8'hc0,8'h80,8'h80,8'hc0,8'h40,8'h80,8'hc0,8'h40,8'hc0,8'h40,8'h80,8'hc0,8'h40,8'h80,8'hc0,8'h40},
	{8'hc0,8'hc0,8'h40,8'h80,8'h80,8'h40,8'hc0,8'h40,8'h80,8'hc0,8'h40,8'h80,8'hc0,8'h40,8'hc0,8'hc0,8'h40,8'hc0,8'h80,8'h40,8'hc0,8'h40,8'h80,8'hc0,8'h40,8'h80,8'h40,8'h40,8'hc0,8'h40,8'h40,8'hc0},
	{8'h40,8'h80,8'hc0,8'h40,8'h80,8'h80,8'h80,8'hc0,8'h40,8'h80,8'hc0,8'h40,8'h80,8'hc0,8'h40,8'h80,8'hc0,8'h40,8'hc0,8'h40,8'h80,8'hc0,8'h40,8'h80,8'hc0,8'h40,8'hc0,8'h40,8'h80,8'hc0,8'h40,8'h40},
	{8'hc0,8'h40,8'hc0,8'hc0,8'h40,8'hc0,8'h80,8'h40,8'hc0,8'h40,8'h80,8'hc0,8'h40,8'h80,8'hc0,8'h40,8'h80,8'hc0,8'h40,8'hc0,8'h40,8'h80,8'hc0,8'h40,8'h80,8'hc0,8'h40,8'hc0,8'h40,8'h40,8'hc0,8'h00},
	{8'h80,8'hc0,8'h40,8'hc0,8'hc0,8'h40,8'hc0,8'h80,8'h80,8'hc0,8'h40,8'h80,8'hc0,8'h40,8'h80,8'hc0,8'h40,8'hc0,8'h80,8'h40,8'hc0,8'h40,8'h80,8'hc0,8'h40,8'h80,8'hc0,8'h40,8'hc0,8'h40,8'h80,8'hc0},
	{8'h40,8'h80,8'hc0,8'h40,8'hc0,8'hc0,8'h40,8'hc0,8'h80,8'h40,8'hc0,8'h40,8'h80,8'hc0,8'h40,8'h80,8'hc0,8'h40,8'hc0,8'hc0,8'h40,8'hc0,8'h40,8'h80,8'hc0,8'h40,8'h80,8'hc0,8'h40,8'hc0,8'h00,8'h40},
	{8'hc0,8'h40,8'h80,8'hc0,8'h40,8'hc0,8'hc0,8'h40,8'hc0,8'h80,8'h80,8'hc0,8'h40,8'h80,8'hc0,8'h40,8'h80,8'hc0,8'h40,8'h80,8'h80,8'h40,8'hc0,8'h40,8'h80,8'hc0,8'h40,8'h80,8'hc0,8'h40,8'hc0,8'h00},
	{8'h80,8'hc0,8'h40,8'h80,8'hc0,8'h40,8'hc0,8'hc0,8'h40,8'hc0,8'h40,8'h40,8'hc0,8'h40,8'h80,8'hc0,8'h40,8'h80,8'hc0,8'h40,8'h80,8'h80,8'h40,8'hc0,8'h40,8'h80,8'hc0,8'h40,8'h80,8'hc0,8'h40,8'hc0},
	{8'h40,8'h80,8'hc0,8'h40,8'h80,8'hc0,8'h40,8'hc0,8'hc0,8'h40,8'hc0,8'h40,8'h80,8'hc0,8'h40,8'h80,8'hc0,8'h40,8'h80,8'hc0,8'h40,8'hc0,8'h80,8'h40,8'hc0,8'h40,8'h80,8'hc0,8'h40,8'h80,8'hc0,8'h40},
	{8'hc0,8'h40,8'h80,8'hc0,8'h40,8'h80,8'hc0,8'h40,8'hc0,8'hc0,8'h40,8'hc0,8'h40,8'h40,8'hc0,8'h40,8'h80,8'hc0,8'h40,8'h80,8'hc0,8'h40,8'hc0,8'h80,8'h40,8'hc0,8'h40,8'h80,8'hc0,8'h40,8'h80,8'hc0},
	{8'h80,8'hc0,8'h00,8'h80,8'hc0,8'h40,8'h80,8'hc0,8'h40,8'hc0,8'hc0,8'h40,8'hc0,8'h40,8'h80,8'hc0,8'h40,8'h80,8'hc0,8'h40,8'h80,8'hc0,8'h40,8'hc0,8'h80,8'h40,8'hc0,8'h40,8'h80,8'hc0,8'h40,8'h80},
	{8'h80,8'h80,8'hc0,8'h40,8'h80,8'hc0,8'h40,8'h80,8'hc0,8'h40,8'hc0,8'hc0,8'h40,8'hc0,8'h40,8'h80,8'hc0,8'h40,8'h80,8'hc0,8'h40,8'h80,8'hc0,8'h40,8'hc0,8'h80,8'h40,8'hc0,8'h00,8'h80,8'hc0,8'h40},
	{8'hc0,8'h80,8'h80,8'hc0,8'h40,8'h80,8'hc0,8'h40,8'h80,8'hc0,8'h40,8'hc0,8'hc0,8'h40,8'hc0,8'h40,8'h80,8'hc0,8'h40,8'h80,8'hc0,8'h40,8'h80,8'hc0,8'h40,8'hc0,8'h40,8'h40,8'hc0,8'h40,8'h80,8'hc0},
	{8'h80,8'hc0,8'h80,8'h80,8'hc0,8'h40,8'h80,8'hc8,8'h40,8'h80,8'hc0,8'h40,8'hc0,8'hc0,8'h40,8'hc0,8'h40,8'h80,8'hc0,8'h40,8'h80,8'hc0,8'h40,8'h80,8'hc0,8'h40,8'hc0,8'h40,8'h80,8'hc0,8'h40,8'h80},
	{8'h80,8'h40,8'hc0,8'h80,8'h80,8'hc0,8'h40,8'h80,8'hc0,8'h40,8'h80,8'hc0,8'h40,8'hc0,8'hc0,8'h40,8'hc0,8'h40,8'h80,8'hc0,8'h40,8'h80,8'hc0,8'h40,8'h80,8'hc0,8'h40,8'hc0,8'h40,8'h80,8'hc0,8'h40}};

 	 
//////////--------------------------------------------------------------------------------------------------------------= 

always_ff@(posedge clk or negedge resetN) 
begin 
	if(!resetN) begin 
		RGBout <=	TRANSPARENT_ENCODING;
	end 
	else begin 
		case (level)
			4'b0001: RGBout <= object_colors[pixelY[4:0]][pixelX[4:0]];          // as it is (red)
			4'b0010: RGBout <= object_colors[pixelY[4:0]][pixelX[4:0]] + 8'h77 ; // blue colors
			4'b0011: RGBout <= object_colors[pixelY[4:0]][pixelX[4:0]] - 8'hA3 ; // green colors
			4'b0000: RGBout <= object_colors[pixelY[4:0]][pixelX[4:0]];          // as it is (red)
		endcase
	end 
end 
 
 
endmodule
