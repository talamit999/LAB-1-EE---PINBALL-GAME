// HartsMatrixBitMap File 
// A two level bitmap. dosplaying harts on the screen FWbruary  2021  
// (c) Technion IIT, Department of Electrical Engineering 2021 



module	StarMatrixBitMap	(	
					input	logic	clk,
					input	logic	resetN,
					input logic	[10:0] offsetX,// offset from top left  position 
					input logic	[10:0] offsetY,
					input	logic	InsideRectangle, //input that the pixel is within a bracket 
					input logic hit,

					output	logic	drawingRequest, //output that the pixel should be dispalyed 
					output	logic	[7:0] RGBout  //rgb value from the bitmap 
 ) ;
 

// Size represented as Number of X and Y bits 
localparam logic [7:0] TRANSPARENT_ENCODING = 8'h00 ;// RGB value in the bitmap representing a transparent pixel 
 /*  end generated by the tool */
 
 localparam logic [7:0] ORANGE = 8'hEC ;
 localparam logic [7:0] PINK = 8'hE2 ;


// the screen is 640*480  or  20 * 15 squares of 32*32  bits ,  we wiil round up to 32*16 and use only the top left 20*15 pixels  
// this is the bitmap  of the maze , if there is a one  the na whole 32*32 rectange will be drawn on the screen 
// all numbers here are hard coded to simplify the  understanding 

logic color_box= 1'b0;//decide the color and change it while collision with ball
							 // 0 -> ORANGE
							 // 1 -> PINK

logic [0:15] [0:15]  MazeBiMapMask= 
{16'b	0000000000000000,
16'b	0000010100000000,
16'b	0000000000000000,
16'b	0000001000000000,
16'b	0000000000000000,
16'b	0000000000000000,
16'b	0000000000000000,
16'b	0000000000000000,
16'b	0000000000000000,
16'b	0000000000000000,
16'b	0000000000000000,
16'b	0000000000000000,
16'b	0000000000000000,
16'b	0000000000000000,
16'b	0000000000000000,
16'b	0000000000000000};


logic[0:31][0:31] object_colors = {
	32'b00000000000000000000000000000000,
	32'b00000000000000000000000000000000,
	32'b00000000000000011000000000000000,
	32'b00000000000000011000000000000000,
	32'b00000000000000111100000000000000,
	32'b00000000000000111100000000000000,
	32'b00000000000001111110000000000000,
	32'b00000000000001111110000000000000,
	32'b00000000000011111111000000000000,
	32'b00000000000011111111000000000000,
	32'b00000000000111111111100000000000,
	32'b00000011111111111111111111000000,
	32'b01111111111111111111111111111110,
	32'b00111111111111111111111111111100,
	32'b00011111111111111111111111111000,
	32'b00001111111111111111111111110000,
	32'b00000111111111111111111111100000,
	32'b00000011111111111111111111000000,
	32'b00000001111111111111111110000000,
	32'b00000000111111111111111100000000,
	32'b00000000111111111111111100000000,
	32'b00000000111111111111111100000000,
	32'b00000000111111111111111100000000,
	32'b00000000111111111111111100000000,
	32'b00000001111111111111111100000000,
	32'b00000001111111111111111110000000,
	32'b00000001111111100111111110000000,
	32'b00000001111110000001111110000000,
	32'b00000001111000000000011110000000,
	32'b00000001100000000000001110000000,
	32'b00000001000000000000000010000000,
	32'b00000000000000000000000000000000};
 

// pipeline (ff) to get the pixel color from the array 	 

//==----------------------------------------------------------------------------------------------------------------=
always_ff@(posedge clk or negedge resetN)
begin
	if(!resetN) begin
		RGBout <= TRANSPARENT_ENCODING;
	end
	else begin
	   // default 
		RGBout <= TRANSPARENT_ENCODING ; 
		
		// change the color if one of the stars hit the ball
		if(hit)
			color_box = ~color_box; 
		
		// only if inside the external bracket and if there is '1' on matrix of stars
		if ((InsideRectangle == 1'b1 ) && (MazeBiMapMask[offsetY[8:5]][offsetX[8:5]] == 1'b1 )) // take bits 5,6,7,8,9,10 from address to select  position in the maze 
			begin
				if(object_colors[offsetY[4:0]][offsetX[4:0]]) begin
					if(color_box)
						RGBout <= PINK;
					else RGBout <= ORANGE;
				end
			end
	end 
end

//==----------------------------------------------------------------------------------------------------------------=
// decide if to draw the pixel or not 
assign drawingRequest = (RGBout != TRANSPARENT_ENCODING ) ? 1'b1 : 1'b0 ;  


endmodule

